* C:\Documents and Settings\All Users\Documents\Softwares\VLSI Softwares\Export dsch2\AdcFlash3bits.sch
* DSCH 2.7a
* created 8/10/2004 3:33:21 PM
*
R1 2 3 50
R2 4 5 50
V1 1 0 DC 1.2
R3 7 4 50
R4 8 7 50
R5 9 8 50
R6 1 6 50
R7 6 9 50
V2 1 0 DC 1.2
R8 5 10 50
*
* Mos models in 0.12�m
* Model 3 n-channel MOS
.MODEL  TN  NMOS
+ LEVEL=3            TPG=+1
+ GAMMA=0.2          THETA=0.5          KAPPA=0.1        ETA=0.002
+ DELTA=0.0          UO=620             VMAX=100E3       VTO=0.35
+ TOX=3e-9           XJ=0.1U            LD=0.00U         NSUB=1E+18
+ NSS=0.2            NFS=7E11
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2
+ CGSO=3.93E-10      CGDO=3.93E-10
* Model 3 p-channel MOS
.MODEL  TP  PMOS
+ LEVEL=3            TPG=-1
+ GAMMA=0.2          THETA=0.5          KAPPA=0.01         ETA=0.001
+ DELTA=0.0          UO=250             VMAX=500E3         VTO=-0.35
+ TOX=3E-9          XJ=0.1U             LD=0.0U             NSUB=1E+18
+ NSS=0.0            NFS=7E11
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
.TRAN 0.1N 50N
* Commands for WinSpice3
* No break in output file
*#set nobreak
* Dump time and volts in "out.txt"
*#print   > out.txt
* Run simulation
*#run
* Show the result in a window
*#plot  
.OPTIONS DELMIN=0 RELTOL=1E-6
.END
